netcdf filter_input {
dimensions:
	member = 50 ;
	metadatalength = 32 ;
	location =  6 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "Field number" ;
		location:dimension = 1 ;
		location:valid_range = 1., 10. ;

	double state(time, member, location) ;
		state:long_name = "the ensemble of model states" ;

	double state_priorinf_mean(time, location) ;
		state_priorinf_mean:long_name = "prior inflation value" ;

	double state_priorinf_sd(time, location) ;
		state_priorinf_sd:long_name = "prior inflation standard deviation" ;

	double state_postinf_mean(time, location) ;
		state_postinf_mean:long_name = "posterior inflation value" ;

	double state_postinf_sd(time, location) ;
		state_postinf_sd:long_name = "posterior inflation standard deviation" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "years" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "none" ;
		advance_to_time:units = "years" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id: $" ;
		:model = "Yasso" ;
		:model_forcing = 8. ;
		:model_deltat = 0.05 ;
		:history = "Varied initial states based on prior drivers" ;
data:

 MemberMetadata =
  "ensemble member       1 ",
  "ensemble member       2 ",
  "ensemble member       3 ",
  "ensemble member       4 ",
  "ensemble member       5 ",
  "ensemble member       6 ",
  "ensemble member       7 ",
  "ensemble member       8 ",
  "ensemble member       9 ",
  "ensemble member       10 ",
  "ensemble member       11 ",
  "ensemble member       12 ",
  "ensemble member       13 ",
  "ensemble member       14 ",
  "ensemble member       15 ",
  "ensemble member       16 ",
  "ensemble member       17 ",
  "ensemble member       18 ",
  "ensemble member       19 ",
  "ensemble member       20 ",
  "ensemble member       21 ",
  "ensemble member       22 ",
  "ensemble member       23 ",
  "ensemble member       24 ",
  "ensemble member       25 ",
  "ensemble member       26 ",
  "ensemble member       27 ",
  "ensemble member       28 ",
  "ensemble member       29 ",
  "ensemble member       30 ",
  "ensemble member       31 ",
  "ensemble member       32 ",
  "ensemble member       33 ",
  "ensemble member       34 ",
  "ensemble member       35 ",
  "ensemble member       36 ",
  "ensemble member       37 ",
  "ensemble member       38 ",
  "ensemble member       39 ",
  "ensemble member       40 ",
  "ensemble member       41 ",
  "ensemble member       42 ",
  "ensemble member       43 ",
  "ensemble member       44 ",
  "ensemble member       45 ",
  "ensemble member       46 ",
  "ensemble member       47 ",
  "ensemble member       48 ",
  "ensemble member       49 ",
  "ensemble member       50 ";

 location = 1, 1, 1, 1, 1, 1 ;

state =
    9.06388820988522, 1.60421823836852, 0.146149008274398, 0.104989565380083, 2.13743961559814, 5.07109178226408, 8.89424077756969, 1.94767818709702, 0.135294070676195, 0.0456684095249975, 2.51939478249638, 4.24620532777511, 12.7790973941131, 1.67029507805282, 0.16198748757122, 0.0900895514407895, 1.84231021530174, 9.01441506174649, 9.79485165216165, 1.18149396833556, 0.156689280387752, 0.0718425441570556, 3.17944243391154, 5.20538342536974, 11.3075662598836, 1.85765192836435, 0.148517612026681, 0.0861537511340312, 2.80502290827492, 6.41022006008358, 9.60495463035634, 1.67142143634031, 0.183225103366211, 0.0936267688636484, 2.15007572029232, 5.50660560149385, 11.2480978573345, 1.49597472505695, 0.146000008249671, 0.11345702203335, 2.94767292618903, 6.54499317580546, 11.4018768373477, 1.51671617519017, 0.197196938753054, 0.146290075727068, 2.87249425453974, 6.66917939313769, 8.60222066527972, 1.42074194072306, 0.202764746499759, 0.0698824053979578, 2.46309084014572, 4.44574073251322, 12.2485991732828, 1.41335333124186, 0.174877757382337, 0.0578149275888591, 3.05717792754558, 7.54537522952421, 7.93824891191587, 0.734932516858013, 0.156785269622457, 0.0696184439867879, 2.72645445392416, 4.25045822752444, 11.5454791644596, 1.26666908952308, 0.112320031737657, 0.125039738140682, 2.58796291347118, 7.45348739158698, 9.49243811442449, 1.29244384154294, 0.142611512702209, 0.0681525169896709, 2.34189361031043, 5.64733663287924, 12.5600828020882, 1.74399035322947, 0.154137624051739, 0.111450316116908, 2.14130192777254, 8.40920258091749, 9.500698765919, 1.63401927064257, 0.190919791934163, 0.0939525056901262, 2.61930609128647, 4.96250110636567, 10.7047805907848, 1.94985422809534, 0.165367348610565, 0.0855507272843109, 1.96644060615545, 6.53756768063913, 7.0043807099513, 1.50957654246381, 0.195856213202089, 0.0803154974609419, 1.23879556745709, 3.97983688936737, 11.7872531550751, 1.29850080809032, 0.127867673172606, 0.091642164255687, 3.34096309548885, 6.92827941406763, 12.5104732624142, 1.7579259347749, 0.186849984252419, 0.102531261507684, 3.59757126162742, 6.8655948202518, 12.0384013131254, 1.95958030651813, 0.207776122662588, 0.104626728746035, 2.16068427056562, 7.60573388463299, 11.2429809299136, 1.56540830711518, 0.218904434773785, 0.0937414755523133, 3.27126702867193, 6.09365968380038, 12.3882912314467, 1.63857634634834, 0.218732653283779, 0.0755664640690684, 3.45189345343927, 7.00352231430622, 11.9107111433516, 1.7980040829446, 0.157110469637356, 0.0885859592211954, 2.1410652947699, 7.72594533677856, 11.0778577385531, 1.88665538050642, 0.180856015754408, 0.073572869857772, 2.26377615492415, 6.67299731751037, 11.4453676548978, 1.6313652806459, 0.160835339689272, 0.10165823227666, 2.22580387997131, 7.32570492231467, 12.8752028392913, 2.10036475095117, 0.181658271128975, 0.0868431796310465, 2.68207315202894, 7.82426348555117, 11.9478157156144, 1.45286744459873, 0.147936181247566, 0.102585409670982, 1.30507096216766, 8.93935571792946, 10.6325942897264, 1.59716016958008, 0.186281838650818, 0.0895956214031869, 2.60826548179101, 6.15129117830129, 11.3519281670974, 1.27108145548767, 0.165949404162416, 0.0738135776771224, 2.60439268068694, 7.23669104908321, 9.26180108254002, 1.88089239779849, 0.110752911163986, 0.0874750713406904, 2.42975305142929, 4.75292765080756, 12.0608583779557, 1.56078021184558, 0.164644738075345, 0.103802654940912, 2.9852569663498, 7.24637380674409, 12.4893694724996, 1.35063730143192, 0.160742321980943, 0.0914960707037578, 2.65173956477344, 8.23475421360957, 11.9347345954297, 1.35408567873394, 0.140951381271657, 0.063413466645745, 2.71761405601402, 7.6586700127643, 11.397852346844, 1.67217005831687, 0.180646359370597, 0.0874769185771283, 2.10626392607225, 7.35129508450713, 11.4061497273988, 1.56758380130359, 0.167995175669632, 0.0769851250132372, 1.8478951782644, 7.74569044714796, 10.3610734993781, 1.72970918677319, 0.160410099819094, 0.0744007158281372, 2.47407554585974, 5.92247795109798, 11.3172491831717, 1.58063576801658, 0.170073380764744, 0.118567661658169, 3.60576505469032, 5.84220731804188, 12.3640467904529, 2.0949701892925, 0.162169605017103, 0.0564210176999792, 2.5487716135656, 7.50171436487773, 10.5416316641642, 1.27806669266472, 0.121758536704557, 0.0904067282757668, 2.17206020902397, 6.87933949749519, 11.2245699084201, 0.862772196482021, 0.163069347752824, 0.0679876296237964, 2.00870351287764, 8.12203722168382, 10.7293357634781, 1.01678025260646, 0.1368570682175, 0.112131529346136, 2.4029307264349, 7.06063618687314, 14.398124773138, 1.79470536433914, 0.158770805482173, 0.11093155051363, 3.41883476939414, 8.91488228340887, 9.98307833184234, 1.83830945408503, 0.152657606418501, 0.107697937570814, 2.38186130832745, 5.50255202544055, 11.5185545283366, 1.41380336289497, 0.153833760547151, 0.11316601719567, 3.286693394603, 6.55105799309581, 8.45862404421457, 1.21250715082431, 0.139607016706969, 0.0899185009528789, 1.92171193382045, 5.09487944190996, 10.4534474382609, 1.72160783579705, 0.16903246342794, 0.114047632670933, 2.16884998186153, 6.27990952450342, 9.0947459220205, 1.64401574381716, 0.166322467441823, 0.111892182880134, 1.76729713091857, 5.40521839696281, 12.4246774896095, 1.373925015324, 0.170564513118138, 0.0498189067381588, 2.09166140322409, 8.73870765120516, 10.8872347173214, 2.00586904212527, 0.18430055443515, 0.088334263934153, 2.93966013264942, 5.66907072417737, 10.3685188003851, 1.19456413983399, 0.106368854462474, 0.0518788621390894, 2.2086571994615, 6.80704974448804 ;

 state_priorinf_mean =
   1, 1, 1, 1, 1, 1 ;

 state_priorinf_sd =
   0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 state_postinf_mean =
   1, 1, 1, 1, 1, 1 ;

 state_postinf_sd =
   0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 time = 1. ;

 advance_to_time = 1. ;
}